<headers>

entity <Name> is

end <Name>;

architecture behave of <Name> is

<component>

<signals>

<stimuli_input>

begin

<clock_gen>

<instance>

<process>

end behave;
